--LIBRARY ieee;
--USE ieee.std_logic_1164.all;
--
--entity contador_Ring is 
--	port
--	(
--		-- Input ports
--		CLK : in std_logic;
--		clr : in STD_LOGIC;
--		EN : IN STD_LOGIC;
--		Putget : in std_logic;
--	
--		-- Output ports
--		Q : out std_logic_vector(2 downto 0)
--	);
--end contador_Ring;
--
--architecture structural of contador_Ring is
--begin
--
--
--
--end structural;